
// Uncomment any testbench for use (by one)


// Counter
//`include "counter-testbench.sv"


// Shift
`include "shift-testbench.sv"


// Shift-get
//`include "shift_gen-testbench.sv"

