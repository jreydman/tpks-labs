
// Uncomment any testbench for use (by one)


// valve [syntax]
//`include "vl-testbench.sv"


// dataflow [syntax]
//`include "df-testbench.sv"


// valve assert test between df and vl modules
//`include "assert-df_vl-testbench.sv"

// mix [syntax]
`include "mix-testbench.sv"
